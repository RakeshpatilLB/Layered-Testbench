`timescale 1ns / 1ps

interface intf(input logic clk, reset);

                
                 logic [31 : 0]  a;
                 logic [31 : 0]  b;
                 logic [31 : 0]  c;
                 logic [31 : 0]  d;

                 logic [31 : 0] a_prim;
                 logic [31 : 0] b_prim;
                 logic [31 : 0] c_prim;
                 logic [31 : 0] d_prim;

endinterface
